--**************************************************************************************--
--					ENSA FES					--
--		             	     Filiere :GSEII					--
--**************************************************************************************--
	-- Title	: bascule D
	-- Project    	: "calculateur de vitesse de rotation d'un moteur"
	-- Block 	: circuit de base
--**************************************************************************************--
	-- File  	: D_BAS.VHD
	-- Authors 	: MIKOU Badr
	-- Created 	: 05/09/2020
--**************************************************************************************--
	-- Description	:
	-- ik ajoute 1 a chaque entrï¿½e.

--**************************************************************************************--


--**************************************************************************************--
--*				     Used Libraries				       *--
--**************************************************************************************--
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;
--**************************************************************************************--
--*				   ENTITY Declaration				       *--
--**************************************************************************************--
ENTITY D_BAS IS PORT (
    rst : IN STD_LOGIC;
    clk : IN STD_LOGIC;
    d   : IN STD_LOGIC;
    q   : OUT STD_LOGIC;
    q_n : OUT STD_LOGIC -- not q
);
END D_BAS;
--**************************************************************************************--
--*				    RTL Description				       *--
--**************************************************************************************--
ARCHITECTURE RTL OF D_BAS IS
BEGIN

    -- le processus de fonctionement 
D_p : PROCESS(CLK)
BEGIN
    IF (rst = '0') THEN
    q   <= '0';
    q_n <= '1'; 
    ELSIF (CLK'EVENT AND CLK = '1') THEN
        q   <= d;
        q_n <= NOT(d);
    END IF;
END PROCESS;

 END RTL;