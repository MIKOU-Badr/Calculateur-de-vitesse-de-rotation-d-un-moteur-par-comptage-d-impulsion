--**************************************************************************************--
--					ENSA FES					--
--		             	     Filiere :GSEII					--
--**************************************************************************************--
	-- Title	: comparateur
	-- Project    	: "calculateur de vitesse de rotation d'un moteur"
    -- Block 	: circuit de base
--**************************************************************************************--
	-- File  	: CMP.VHD
	-- Authors 	: MIKOU Badr
	-- Created 	: 04/09/2020
--**************************************************************************************--
	-- Description	:
	-- la sortie y prend 1 si in0 = in1.
	-- 
	 
--**************************************************************************************--


--**************************************************************************************--
--*				     Used Libraries				       *--
--**************************************************************************************--
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;
--**************************************************************************************--
--*				   ENTITY Declaration				       *--
--**************************************************************************************--

ENTITY CMP IS PORT (
	in0 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
	in1 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
	y   : OUT STD_LOGIC);
END CMP;

--**************************************************************************************--
--*				    RTL Description				       *--
--**************************************************************************************--

ARCHITECTURE RTL OF CMP IS
BEGIN

y <= '1' WHEN (in1 = in0) ELSE
     '0';
     
 END RTL;