--**************************************************************************************--
--					ENSA FES					--
--		             	     Filiere :GSEII					--
--**************************************************************************************--
	-- Title	: aditionneur de 1
	-- Project    	: "calculateur de vitesse de rotation d'un moteur"
	-- Block 	: circuit de base
--**************************************************************************************--
	-- File  	: ADD_1_GEN.VHD
	-- Authors 	: MIKOU Badr
	-- Created 	: 04/09/2020
--**************************************************************************************--
	-- Description	:
	-- ik ajoute 1 a chaque entr�e.

--**************************************************************************************--


--**************************************************************************************--
--*				     Used Libraries				       *--
--**************************************************************************************--
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;
--**************************************************************************************--
--*				   ENTITY Declaration				       *--
--**************************************************************************************--
ENTITY ADD_1_GEN IS GENERIC ( 
	n : INTEGER := 5
);
PORT (
    a : IN STD_LOGIC_VECTOR(n-1 DOWNTO 0);
	s : OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0)
);
END ADD_1_GEN;
--**************************************************************************************--
--*				    RTL Description				       *--
--**************************************************************************************--
ARCHITECTURE RTL OF ADD_1_GEN IS
    
    SIGNAL sig_1 :STD_LOGIC_VECTOR(n-1 DOWNTO 0);
    
    BEGIN
        sig_1 <= a + '1';
        s <= sig_1;
 END RTL;